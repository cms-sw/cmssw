-- alp2,alp1,name,tl2,h2,h1,bl1,tl1,bl2,phi,dz,theta
