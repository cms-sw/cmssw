-- name,dx2,dx1,dy1,dz,dy2
