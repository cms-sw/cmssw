-- dz,name,dx,dy
