-- deltaPhi,name,numSide,startPhi,RZ_or_ZS
