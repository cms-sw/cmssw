-- sequence_no,rMin,z,rMax,polycone_solid_name,polyhedra_solid_name
