-- deltaPhi,name,startPhi,RZ_or_ZS
