-- name,rMin1,rMax1,rMax2,dz,deltaPhi,startPhi,rMin2
