-- name,operation,solidA,solidB,x,y,z,ro
