-- dz,name,dx,dy
