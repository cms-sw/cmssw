-- rMin,name,rMax,deltaPhi,dz,startPhi
